----------------------------------------------------------------------------------
-- Company: UTCN
-- Engineer: Raluca Adam
-- 
-- Create Date: 05/03/2024 04:29:22 PM
-- Design Name: Flags Register
-- Module Name: FlagsRegister - Behavioral
-- Project Name: Microcontroller
-- Target Devices: Artix-7 100T
-- Tool Versions: 
-- Description: 
--          register stores the ZERO and CARRY flags generated by the ALU
--          asynhrounous RESET
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity FlagsRegister is
    Port ( ZFIN : in STD_LOGIC;
           CFIN : in STD_LOGIC;
           ZFOUT : out STD_LOGIC;
           CFOUT : out STD_LOGIC;
           CLK : in STD_LOGIC;
           RESET : in STD_LOGIC);
end FlagsRegister;

architecture Behavioral of FlagsRegister is

begin
    process(CLK, RESET)
    variable zero, carry: std_logic := '0';
    begin
        if RESET = '1' then 
            zero := '0';
            carry := '0';
        else
            if (CLK'event) and (CLK = '1') then
                zero := ZFIN;
                carry := CFIN;
            end if;
        end if;
        ZFOUT <= zero;
        CFOUT <= carry;
    end process;
end Behavioral;